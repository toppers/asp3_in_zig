/*
 *		テスト用プラットフォーム（カーネルの整合性検査付き）のコンポー
 *		ネント記述ファイル
 *
 *  $Id: test_pf_bitkernel.cdl 882 2018-02-01 09:55:37Z ertl-hiro $
 */

/*
 *  テスト用プラットフォームのコンポーネント記述ファイル
 */
import("test_pf.cdl");

/*
 *  カーネルの整合性検査のセルタイプと組上げ記述
 */
[singleton]
celltype tBitKernel {
	entry	sBuiltInTest	eBuiltInTest;
};

cell tBitKernel BitKernel {
	eBuiltInTest <= TestService.cBuiltInTest;	/* テストサービスに接続 */
};
